`default_nettype none

// start your project from here.
module top (
    input wire 
);



endmodule
